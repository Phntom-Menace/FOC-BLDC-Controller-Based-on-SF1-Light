// Verilog netlist created by Tang Dynasty v5.6.71036
// Fri Nov 10 01:09:53 2023

`timescale 1ns / 1ps
module Divider
  (
  clk,
  denominator,
  numerator,
  rst,
  start,
  done,
  quotient,
  remainder
  );

  input clk;
  input [5:0] denominator;
  input [17:0] numerator;
  input rst;
  input start;
  output done;
  output [17:0] quotient;
  output [5:0] remainder;

  parameter S_DEN = "UNSIGNED";
  parameter S_NUM = "UNSIGNED";
  parameter W_DEN = 6;
  parameter W_NUM = 18;
  // localparam W_CNT = 5;
  wire [4:0] al_1deac949;
  wire [4:0] al_d0dc52fd;
  wire [22:0] al_11033702;
  wire [22:0] al_1c1b24e7;
  wire [17:0] al_1315ed94;
  wire [17:0] al_9bfb1470;
  wire [22:0] al_c67bebad;
  wire [17:0] al_327525b3;
  wire al_9673d977;
  wire al_a9fbe072;
  wire al_3973d008;
  wire al_4c40b6e5;
  wire al_d63e42fe;
  wire al_b4fc1000;
  wire al_ab829401;
  wire al_b7ca2ed;
  wire al_22a7ce9f;
  wire al_f5902502;
  wire al_b83a67b2;
  wire al_540b209;
  wire al_27e1f3bc;
  wire al_e64e5f1c;
  wire al_e761a920;
  wire al_42ead886;
  wire al_f5a327ab;
  wire al_b23e28b5;
  wire al_283f8d98;
  wire al_516747bd;
  wire al_88a2e01;
  wire al_424d2e3a;
  wire al_5d3a435a;
  wire al_4a5ad68f;
  wire al_76de0dc5;
  wire al_8d09201;
  wire al_373410a0;
  wire al_34afb8ef;
  wire al_cba3eae;
  wire al_778bfe34;
  wire al_7f34b742;
  wire al_dd7c9c08;
  wire al_6b6ab26e;
  wire al_4331c4e0;
  wire al_a5be61f4;
  wire al_f577d7c;
  wire al_f39a7e9;
  wire al_9762a925;
  wire al_ef2ad0c3;
  wire al_e7f7dbb1;
  wire al_b1f223c3;
  wire al_e7086bfe;
  wire al_114eba31;
  wire al_c61b4192;
  wire al_82473adc;
  wire al_b5f6bee4;

  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    al_dc50342 (
    .a(al_82473adc),
    .b(al_1deac949[2]),
    .c(al_1deac949[3]),
    .d(al_1deac949[4]),
    .o(al_114eba31));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_f17cd423 (
    .a(al_1deac949[2]),
    .b(al_1deac949[3]),
    .o(al_b5f6bee4));
  AL_MAP_LUT5 #(
    .EQN("~(~B*~(~C*~(~E*~D*A)))"),
    .INIT(32'hcfcfcfcd))
    al_b4279277 (
    .a(al_b5f6bee4),
    .b(start),
    .c(al_1deac949[0]),
    .d(al_1deac949[1]),
    .e(al_1deac949[4]),
    .o(al_d0dc52fd[0]));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    al_147e6a1b (
    .a(start),
    .b(al_1deac949[0]),
    .c(al_1deac949[1]),
    .o(al_d0dc52fd[1]));
  AL_MAP_LUT5 #(
    .EQN("(~B*(A*~(C)*~((E*~D))+~(A)*C*~((E*~D))+~(A)*C*(E*~D)))"),
    .INIT(32'h12101212))
    al_c8620855 (
    .a(al_82473adc),
    .b(start),
    .c(al_1deac949[2]),
    .d(al_1deac949[3]),
    .e(al_1deac949[4]),
    .o(al_d0dc52fd[2]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    al_6614de08 (
    .a(al_82473adc),
    .b(start),
    .c(al_1deac949[2]),
    .d(al_1deac949[3]),
    .o(al_d0dc52fd[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_6dc5f615 (
    .a(al_1deac949[0]),
    .b(al_1deac949[1]),
    .o(al_82473adc));
  AL_MAP_LUT5 #(
    .EQN("(~B*(A*C*D*~(E)+~(A)*~(C)*~(D)*E+~(A)*C*~(D)*E+A*C*~(D)*E+~(A)*~(C)*D*E+A*~(C)*D*E+~(A)*C*D*E))"),
    .INIT(32'h13312000))
    al_4a3f31d6 (
    .a(al_82473adc),
    .b(start),
    .c(al_1deac949[2]),
    .d(al_1deac949[3]),
    .e(al_1deac949[4]),
    .o(al_d0dc52fd[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_d2344c96 (
    .a(denominator[0]),
    .b(start),
    .c(al_11033702[18]),
    .o(al_1c1b24e7[17]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_faf89982 (
    .a(denominator[1]),
    .b(start),
    .c(al_11033702[19]),
    .o(al_1c1b24e7[18]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_22b9e4c0 (
    .a(denominator[2]),
    .b(start),
    .c(al_11033702[20]),
    .o(al_1c1b24e7[19]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_b1b9ffd0 (
    .a(denominator[3]),
    .b(start),
    .c(al_11033702[21]),
    .o(al_1c1b24e7[20]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_b2cd7517 (
    .a(denominator[4]),
    .b(start),
    .c(al_11033702[22]),
    .o(al_1c1b24e7[21]));
  AL_DFF_0 al_35b11324 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_114eba31),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(done));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    al_2c0796e5 (
    .a(1'b1),
    .o({al_9673d977,open_n2}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_c203f32c (
    .a(al_11033702[4]),
    .b(al_1315ed94[4]),
    .c(al_d63e42fe),
    .o({al_b4fc1000,open_n3}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_5a2e66a8 (
    .a(al_11033702[5]),
    .b(al_1315ed94[5]),
    .c(al_b4fc1000),
    .o({al_ab829401,open_n4}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_2f287d12 (
    .a(al_11033702[6]),
    .b(al_1315ed94[6]),
    .c(al_ab829401),
    .o({al_b7ca2ed,open_n5}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_9ce86edd (
    .a(al_11033702[7]),
    .b(al_1315ed94[7]),
    .c(al_b7ca2ed),
    .o({al_22a7ce9f,open_n6}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_29f6525 (
    .a(al_11033702[8]),
    .b(al_1315ed94[8]),
    .c(al_22a7ce9f),
    .o({al_f5902502,open_n7}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_f171b4f4 (
    .a(al_11033702[0]),
    .b(al_1315ed94[0]),
    .c(al_9673d977),
    .o({al_a9fbe072,open_n8}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e9c7012b (
    .a(al_11033702[9]),
    .b(al_1315ed94[9]),
    .c(al_f5902502),
    .o({al_b83a67b2,open_n9}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_4226b3d1 (
    .a(al_11033702[10]),
    .b(al_1315ed94[10]),
    .c(al_b83a67b2),
    .o({al_540b209,open_n10}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_3f6fc47e (
    .a(al_11033702[11]),
    .b(al_1315ed94[11]),
    .c(al_540b209),
    .o({al_27e1f3bc,open_n11}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e17073e0 (
    .a(al_11033702[12]),
    .b(al_1315ed94[12]),
    .c(al_27e1f3bc),
    .o({al_e64e5f1c,open_n12}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_ba5a9770 (
    .a(al_11033702[13]),
    .b(al_1315ed94[13]),
    .c(al_e64e5f1c),
    .o({al_e761a920,open_n13}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_cb976531 (
    .a(al_11033702[14]),
    .b(al_1315ed94[14]),
    .c(al_e761a920),
    .o({al_42ead886,open_n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e5cd5640 (
    .a(al_11033702[15]),
    .b(al_1315ed94[15]),
    .c(al_42ead886),
    .o({al_f5a327ab,open_n15}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e4d1cd55 (
    .a(al_11033702[16]),
    .b(al_1315ed94[16]),
    .c(al_f5a327ab),
    .o({al_b23e28b5,open_n16}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_dc7e8c2c (
    .a(al_11033702[17]),
    .b(al_1315ed94[17]),
    .c(al_b23e28b5),
    .o({al_283f8d98,open_n17}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_9ed345ca (
    .a(al_11033702[18]),
    .b(1'b0),
    .c(al_283f8d98),
    .o({al_516747bd,open_n18}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_441ad9b2 (
    .a(al_11033702[1]),
    .b(al_1315ed94[1]),
    .c(al_a9fbe072),
    .o({al_3973d008,open_n19}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_36cc28eb (
    .a(al_11033702[19]),
    .b(1'b0),
    .c(al_516747bd),
    .o({al_88a2e01,open_n20}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_e18ee10 (
    .a(al_11033702[20]),
    .b(1'b0),
    .c(al_88a2e01),
    .o({al_424d2e3a,open_n21}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_99bd7325 (
    .a(al_11033702[21]),
    .b(1'b0),
    .c(al_424d2e3a),
    .o({al_5d3a435a,open_n22}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_8aa83152 (
    .a(al_11033702[22]),
    .b(1'b0),
    .c(al_5d3a435a),
    .o({al_4a5ad68f,open_n23}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_1c94cea5 (
    .a(1'b0),
    .b(1'b1),
    .c(al_4a5ad68f),
    .o({open_n24,al_c61b4192}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_9395428b (
    .a(al_11033702[2]),
    .b(al_1315ed94[2]),
    .c(al_3973d008),
    .o({al_4c40b6e5,open_n25}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    al_f7ac689a (
    .a(al_11033702[3]),
    .b(al_1315ed94[3]),
    .c(al_4c40b6e5),
    .o({al_d63e42fe,open_n26}));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_affc23c8 (
    .a(numerator[0]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[0]),
    .e(al_c67bebad[0]),
    .o(al_9bfb1470[0]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_7e4247d5 (
    .a(numerator[10]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[10]),
    .e(al_c67bebad[10]),
    .o(al_9bfb1470[10]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_8f76e334 (
    .a(numerator[11]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[11]),
    .e(al_c67bebad[11]),
    .o(al_9bfb1470[11]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_43c29c9e (
    .a(numerator[12]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[12]),
    .e(al_c67bebad[12]),
    .o(al_9bfb1470[12]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_dcb75b0 (
    .a(numerator[13]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[13]),
    .e(al_c67bebad[13]),
    .o(al_9bfb1470[13]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_e1773c9b (
    .a(numerator[14]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[14]),
    .e(al_c67bebad[14]),
    .o(al_9bfb1470[14]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_8e3693cb (
    .a(numerator[15]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[15]),
    .e(al_c67bebad[15]),
    .o(al_9bfb1470[15]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_79948be9 (
    .a(numerator[16]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[16]),
    .e(al_c67bebad[16]),
    .o(al_9bfb1470[16]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_cd0015f2 (
    .a(numerator[17]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[17]),
    .e(al_c67bebad[17]),
    .o(al_9bfb1470[17]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_db832082 (
    .a(numerator[1]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[1]),
    .e(al_c67bebad[1]),
    .o(al_9bfb1470[1]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_3e04c0e7 (
    .a(numerator[2]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[2]),
    .e(al_c67bebad[2]),
    .o(al_9bfb1470[2]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_b86e3fac (
    .a(numerator[3]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[3]),
    .e(al_c67bebad[3]),
    .o(al_9bfb1470[3]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_1f499def (
    .a(numerator[4]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[4]),
    .e(al_c67bebad[4]),
    .o(al_9bfb1470[4]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_8f1711f3 (
    .a(numerator[5]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[5]),
    .e(al_c67bebad[5]),
    .o(al_9bfb1470[5]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_6e1c653d (
    .a(numerator[6]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[6]),
    .e(al_c67bebad[6]),
    .o(al_9bfb1470[6]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_b46e3fd7 (
    .a(numerator[7]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[7]),
    .e(al_c67bebad[7]),
    .o(al_9bfb1470[7]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_d21f8608 (
    .a(numerator[8]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[8]),
    .e(al_c67bebad[8]),
    .o(al_9bfb1470[8]));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'hbbb88b88))
    al_42e41119 (
    .a(numerator[9]),
    .b(start),
    .c(al_c61b4192),
    .d(al_1315ed94[9]),
    .e(al_c67bebad[9]),
    .o(al_9bfb1470[9]));
  AL_DFF_0 al_b26d62bf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[0]));
  AL_DFF_0 al_809f7104 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[1]));
  AL_DFF_0 al_c1468025 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[2]));
  AL_DFF_0 al_c19d8344 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[3]));
  AL_DFF_0 al_ca1eda73 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_d0dc52fd[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1deac949[4]));
  AL_DFF_0 al_b40e8e05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[9]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[8]));
  AL_DFF_0 al_2259e8d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[10]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[9]));
  AL_DFF_0 al_5f624aaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[11]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[10]));
  AL_DFF_0 al_d532b054 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[12]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[11]));
  AL_DFF_0 al_9d987fc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[13]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[12]));
  AL_DFF_0 al_220744cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[14]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[13]));
  AL_DFF_0 al_e241f44a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[15]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[14]));
  AL_DFF_0 al_897da5eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[16]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[15]));
  AL_DFF_0 al_9e863954 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[17]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[16]));
  AL_DFF_0 al_a186fcad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[17]));
  AL_DFF_0 al_fd544ba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[1]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[0]));
  AL_DFF_0 al_21ba363c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[18]));
  AL_DFF_0 al_c602bc36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[19]));
  AL_DFF_0 al_be443a52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[20]));
  AL_DFF_0 al_961a8bb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c1b24e7[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_11033702[21]));
  AL_DFF_0 al_6d594c9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[5]),
    .en(1'b1),
    .sr(~start),
    .ss(1'b0),
    .q(al_11033702[22]));
  AL_DFF_0 al_40ebe0d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[2]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[1]));
  AL_DFF_0 al_b4cd3408 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[3]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[2]));
  AL_DFF_0 al_16607eff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[4]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[3]));
  AL_DFF_0 al_2e1082f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[5]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[4]));
  AL_DFF_0 al_806f02ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[6]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[5]));
  AL_DFF_0 al_e97bb64b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[7]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[6]));
  AL_DFF_0 al_f7f2da08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11033702[8]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_11033702[7]));
  AL_DFF_0 al_596b0fc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[8]));
  AL_DFF_0 al_5cfa2c1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[9]));
  AL_DFF_0 al_c56c02f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[10]));
  AL_DFF_0 al_60ec2662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[11]));
  AL_DFF_0 al_ea3f598e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[12]));
  AL_DFF_0 al_dd4ae85d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[13]));
  AL_DFF_0 al_e2aa8055 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[14]));
  AL_DFF_0 al_82aa8ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[15]));
  AL_DFF_0 al_7f911c70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[16]));
  AL_DFF_0 al_8908ba38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[17]));
  AL_DFF_0 al_16ad90bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[0]));
  AL_DFF_0 al_e1044ec0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[1]));
  AL_DFF_0 al_16da6de4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[2]));
  AL_DFF_0 al_e819e904 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[3]));
  AL_DFF_0 al_4990808d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[4]));
  AL_DFF_0 al_d51e17ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[5]));
  AL_DFF_0 al_b67f884b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[6]));
  AL_DFF_0 al_ff3308ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9bfb1470[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1315ed94[7]));
  AL_DFF_0 al_c1e3ea45 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[8]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[8]));
  AL_DFF_0 al_b7aa029f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[9]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[9]));
  AL_DFF_0 al_2f4f18cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[10]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[10]));
  AL_DFF_0 al_42a7eb97 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[11]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[11]));
  AL_DFF_0 al_f77c099a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[12]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[12]));
  AL_DFF_0 al_6893ba8f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[13]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[13]));
  AL_DFF_0 al_d6d1e991 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[14]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[14]));
  AL_DFF_0 al_4d3bf6cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[15]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[15]));
  AL_DFF_0 al_aa8c310 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[16]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[16]));
  AL_DFF_0 al_d8095998 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[17]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[17]));
  AL_DFF_0 al_53efe64b (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[0]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[0]));
  AL_DFF_0 al_26890f76 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[1]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[1]));
  AL_DFF_0 al_802c7023 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[2]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[2]));
  AL_DFF_0 al_9c45670 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[3]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[3]));
  AL_DFF_0 al_b0a0e999 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[4]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[4]));
  AL_DFF_0 al_739d9f2f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[5]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[5]));
  AL_DFF_0 al_7f9eee7d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[6]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[6]));
  AL_DFF_0 al_741313a7 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[7]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[7]));
  AL_DFF_0 al_ce6e5997 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[7]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[8]));
  AL_DFF_0 al_7c322425 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[8]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[9]));
  AL_DFF_0 al_1f65ec13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[9]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[10]));
  AL_DFF_0 al_63457b5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[10]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[11]));
  AL_DFF_0 al_11fe6cd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[11]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[12]));
  AL_DFF_0 al_9cfb6f54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[12]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[13]));
  AL_DFF_0 al_40b705d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[13]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[14]));
  AL_DFF_0 al_cbb21b57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[14]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[15]));
  AL_DFF_0 al_a743530c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[15]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[16]));
  AL_DFF_0 al_50032887 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[16]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[17]));
  AL_DFF_0 al_5e904a35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c61b4192),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[0]));
  AL_DFF_0 al_116f1db3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[0]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[1]));
  AL_DFF_0 al_6c993e82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[1]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[2]));
  AL_DFF_0 al_23963ea6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[2]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[3]));
  AL_DFF_0 al_6c25cf29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[3]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[4]));
  AL_DFF_0 al_e7cc423c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[4]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[5]));
  AL_DFF_0 al_2c6ea385 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[5]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[6]));
  AL_DFF_0 al_a356779f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_327525b3[6]),
    .en(1'b1),
    .sr(start),
    .ss(1'b0),
    .q(al_327525b3[7]));
  AL_DFF_0 al_cbbb4490 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[0]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[0]));
  AL_DFF_0 al_30153836 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[1]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[1]));
  AL_DFF_0 al_37ead40d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[2]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[2]));
  AL_DFF_0 al_7625712c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[3]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[3]));
  AL_DFF_0 al_2531de5d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[4]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[4]));
  AL_DFF_0 al_2ccbdc6d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_1315ed94[5]),
    .en(al_114eba31),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[5]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8b9c8457 (
    .a(al_1315ed94[7]),
    .b(al_11033702[7]),
    .c(al_dd7c9c08),
    .o({al_6b6ab26e,al_c67bebad[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5e613dd7 (
    .a(al_1315ed94[8]),
    .b(al_11033702[8]),
    .c(al_6b6ab26e),
    .o({al_4331c4e0,al_c67bebad[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_27c8842d (
    .a(al_1315ed94[9]),
    .b(al_11033702[9]),
    .c(al_4331c4e0),
    .o({al_a5be61f4,al_c67bebad[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_462a01f1 (
    .a(al_1315ed94[10]),
    .b(al_11033702[10]),
    .c(al_a5be61f4),
    .o({al_f577d7c,al_c67bebad[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9b3bce39 (
    .a(al_1315ed94[11]),
    .b(al_11033702[11]),
    .c(al_f577d7c),
    .o({al_f39a7e9,al_c67bebad[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f829bb24 (
    .a(al_1315ed94[12]),
    .b(al_11033702[12]),
    .c(al_f39a7e9),
    .o({al_9762a925,al_c67bebad[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cc29264d (
    .a(al_1315ed94[13]),
    .b(al_11033702[13]),
    .c(al_9762a925),
    .o({al_ef2ad0c3,al_c67bebad[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ee4a1d93 (
    .a(al_1315ed94[14]),
    .b(al_11033702[14]),
    .c(al_ef2ad0c3),
    .o({al_e7f7dbb1,al_c67bebad[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_154312aa (
    .a(al_1315ed94[15]),
    .b(al_11033702[15]),
    .c(al_e7f7dbb1),
    .o({al_b1f223c3,al_c67bebad[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17566e78 (
    .a(al_1315ed94[16]),
    .b(al_11033702[16]),
    .c(al_b1f223c3),
    .o({al_e7086bfe,al_c67bebad[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_f5224f5b (
    .a(1'b0),
    .o({al_76de0dc5,open_n29}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_38657e34 (
    .a(al_1315ed94[17]),
    .b(al_11033702[17]),
    .c(al_e7086bfe),
    .o({open_n30,al_c67bebad[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e6e3dfcf (
    .a(al_1315ed94[0]),
    .b(al_11033702[0]),
    .c(al_76de0dc5),
    .o({al_8d09201,al_c67bebad[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_68abff86 (
    .a(al_1315ed94[1]),
    .b(al_11033702[1]),
    .c(al_8d09201),
    .o({al_373410a0,al_c67bebad[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8de058bd (
    .a(al_1315ed94[2]),
    .b(al_11033702[2]),
    .c(al_373410a0),
    .o({al_34afb8ef,al_c67bebad[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bbd4c846 (
    .a(al_1315ed94[3]),
    .b(al_11033702[3]),
    .c(al_34afb8ef),
    .o({al_cba3eae,al_c67bebad[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_222b6767 (
    .a(al_1315ed94[4]),
    .b(al_11033702[4]),
    .c(al_cba3eae),
    .o({al_778bfe34,al_c67bebad[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9c7fbfa5 (
    .a(al_1315ed94[5]),
    .b(al_11033702[5]),
    .c(al_778bfe34),
    .o({al_7f34b742,al_c67bebad[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fd218d47 (
    .a(al_1315ed94[6]),
    .b(al_11033702[6]),
    .c(al_7f34b742),
    .o({al_dd7c9c08,al_c67bebad[6]}));

endmodule 

